    Mac OS X            	   2  �     �                                    ATTR     �   �   K                  �   ;  com.apple.quarantine    �     com.apple.lastuseddate#PS 44E0081;61b16cd6;WhatsApp;246A38F1-56F2-44E9-8DC0-132B60F1FB7A�J�a    +T                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         This resource fork intentionally left blank                                                                                                                                                                                                                            ��